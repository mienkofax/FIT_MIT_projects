
//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_in_wire_en_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_wire_en_v1 (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output [width-1:0] d;
  output             lz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;

endmodule


//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_in_wire_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_in_wire_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule


//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_out_stdreg_en_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_stdreg_en_v1 (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  input  [width-1:0] d;
  output             lz;
  output [width-1:0] z;

  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;

endmodule



//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Block 1R1W Read Before Write RAM with common clock
module BLOCK_1R1W_RBW
#(
parameter data_width = 8,
parameter addr_width = 7,
parameter depth = 128
)(
	radr, wadr, d, we, re, clk, q
);

	input [addr_width-1:0] radr;
	input [addr_width-1:0] wadr;
	input [data_width-1:0] d;
	input we;
	input re;
	input clk;
	output[data_width-1:0] q;

	reg [data_width-1:0] q;

	(* ram_style = "block" *)
	reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block_ram"
	//pragma attribute mem block_ram true
		
	always @(posedge clk) begin
		if (we) begin
			mem[wadr] <= d; // Write port
		end
		if (re) begin
			q <= mem[radr] ; // read port
		end
	end

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0c/745553 Production Release
//  HLS Date:       Wed Oct 11 16:38:17 PDT 2017
// 
//  Generated by:   Fitkit@DESKTOP-NJUNEBJ
//  Generated date: Tue Dec 19 09:42:46 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_10_640_7_gen
// ------------------------------------------------------------------


module Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_10_640_7_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [2:0] d;
  output [9:0] wadr;
  output re;
  input [2:0] q;
  output [9:0] radr;
  input [9:0] radr_d;
  input [9:0] wadr_d;
  input [2:0] d_d;
  input we_d;
  input re_d;
  output [2:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_32_9_512_4_gen
// ------------------------------------------------------------------


module Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_32_9_512_4_gen (
  we, d, q, adr, adr_d, d_d, we_d, q_d, ram_rw_A_internal_RMASK_B_d
);
  output we;
  output [31:0] d;
  input [31:0] q;
  output [8:0] adr;
  input [8:0] adr_d;
  input [31:0] d_d;
  input we_d;
  output [31:0] q_d;
  input ram_rw_A_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign q_d = q;
  assign adr = (adr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    filter_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module filter_core_core_fsm (
  clk, rst, fsm_output, buffer_buf_vinit_C_1_tr0
);
  input clk;
  input rst;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;
  input buffer_buf_vinit_C_1_tr0;


  // FSM State Type Declaration for filter_core_core_fsm_1
  parameter
    core_rlp_C_0 = 3'd0,
    buffer_buf_vinit_C_0 = 3'd1,
    buffer_buf_vinit_C_1 = 3'd2,
    main_C_0 = 3'd3,
    main_C_1 = 3'd4,
    main_C_2 = 3'd5,
    main_C_3 = 3'd6;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : filter_core_core_fsm_1
    case (state_var)
      buffer_buf_vinit_C_0 : begin
        fsm_output = 7'b10;
        state_var_NS = buffer_buf_vinit_C_1;
      end
      buffer_buf_vinit_C_1 : begin
        fsm_output = 7'b100;
        if ( buffer_buf_vinit_C_1_tr0 ) begin
          state_var_NS = buffer_buf_vinit_C_0;
        end
        else begin
          state_var_NS = main_C_0;
        end
      end
      main_C_0 : begin
        fsm_output = 7'b1000;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 7'b10000;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 7'b100000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 7'b1000000;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 7'b1;
        state_var_NS = buffer_buf_vinit_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    filter_core
// ------------------------------------------------------------------


module filter_core (
  clk, rst, in_data_rsc_z, in_data_rsc_lz, in_data_vld_rsc_z, out_data_rsc_z, out_data_rsc_lz,
      mcu_data_rsci_adr_d, mcu_data_rsci_d_d, mcu_data_rsci_we_d, mcu_data_rsci_q_d,
      mcu_data_rsci_ram_rw_A_internal_RMASK_B_d, buffer_buf_rsci_radr_d, buffer_buf_rsci_wadr_d,
      buffer_buf_rsci_d_d, buffer_buf_rsci_we_d, buffer_buf_rsci_re_d, buffer_buf_rsci_q_d
);
  input clk;
  input rst;
  input [2:0] in_data_rsc_z;
  output in_data_rsc_lz;
  input in_data_vld_rsc_z;
  output [2:0] out_data_rsc_z;
  output out_data_rsc_lz;
  output [8:0] mcu_data_rsci_adr_d;
  output [31:0] mcu_data_rsci_d_d;
  output mcu_data_rsci_we_d;
  input [31:0] mcu_data_rsci_q_d;
  output mcu_data_rsci_ram_rw_A_internal_RMASK_B_d;
  output [9:0] buffer_buf_rsci_radr_d;
  output [9:0] buffer_buf_rsci_wadr_d;
  output [2:0] buffer_buf_rsci_d_d;
  output buffer_buf_rsci_we_d;
  output buffer_buf_rsci_re_d;
  input [2:0] buffer_buf_rsci_q_d;


  // Interconnect Declarations
  reg in_data_rsci_ld;
  wire [2:0] in_data_rsci_d;
  wire in_data_vld_rsci_d;
  reg out_data_rsci_ld;
  reg out_data_rsci_d_0;
  wire [6:0] fsm_output;
  wire if_if_if_and_tmp;
  wire [2:0] pixel_processing_mod10_acc_3_tmp;
  wire [3:0] nl_pixel_processing_mod10_acc_3_tmp;
  wire and_tmp;
  wire or_dcpl_1;
  wire and_dcpl_41;
  wire or_dcpl_54;
  wire nor_tmp_5;
  wire nor_tmp_6;
  wire mux_tmp_6;
  wire or_dcpl_75;
  wire or_dcpl_80;
  wire or_dcpl_81;
  wire or_dcpl_87;
  wire and_dcpl_101;
  wire or_dcpl_124;
  wire and_dcpl_126;
  wire or_tmp_35;
  wire or_tmp_49;
  reg mcu_ready_sva;
  reg [2:0] pixel_processing_threshold_sva;
  reg [31:0] pixel_processing_frame_sva;
  wire [32:0] nl_pixel_processing_frame_sva;
  reg [8:0] system_input_c_sva;
  reg [8:0] system_input_c_filter_sva;
  reg [7:0] system_input_r_sva;
  reg [7:0] system_input_r_filter_sva;
  reg system_input_output_vld_sva;
  reg [2:0] system_input_window_4_sva;
  reg [2:0] system_input_window_3_sva;
  reg [2:0] system_input_window_5_sva;
  reg [2:0] system_input_window_6_sva;
  reg [2:0] system_input_window_7_sva;
  reg [2:0] system_input_window_8_sva;
  reg [9:0] buffer_buf_vinit_ndx_sva;
  reg buffer_sel_1_sva;
  reg else_io_read_in_data_vld_rsc_svs;
  reg [2:0] system_input_din_sva_1;
  reg buffer_sel_1_sva_dfm;
  reg [2:0] buffer_t0_sva_1;
  reg clip_window_ac_int_cctor_2_sva_1;
  reg clip_window_clip_window_and_1_cse_sva_1;
  reg clip_window_unequal_tmp_2;
  reg system_input_output_vld_sva_dfm;
  reg system_input_land_1_lpi_1_dfm_1;
  reg [2:0] median_max2_5_1_lpi_1_dfm;
  reg [2:0] median_max_4_2_lpi_1_dfm;
  reg [2:0] median_max2_3_2_lpi_1_dfm;
  reg [2:0] median_max_2_2_lpi_1_dfm;
  reg [2:0] median_max2_1_lpi_1_dfm;
  reg [2:0] median_max_4_1_lpi_1_dfm;
  reg [2:0] median_max_6_lpi_1_dfm;
  reg [2:0] median_max_5_3_lpi_1_dfm;
  reg [2:0] median_max_7_lpi_1_dfm;
  reg pixel_processing_if_2_land_lpi_1_dfm_1;
  reg buffer_buf_buffer_buf_nor_itm_1;
  reg [9:0] buffer_buf_acc_itm_2;
  wire [10:0] nl_buffer_buf_acc_itm_2;
  reg [2:0] median_max_5_lpi_1_dfm_5;
  reg asn_itm;
  reg else_io_read_in_data_vld_rsc_svs_st_1;
  reg [3:0] buffer_acc_1_itm_2;
  wire [4:0] nl_buffer_acc_1_itm_2;
  reg [3:0] buffer_acc_3_itm_2;
  wire [4:0] nl_buffer_acc_3_itm_2;
  reg [5:0] buffer_slc_buffer_c_5_0_1_itm_2;
  reg system_input_output_vld_sva_dfm_st_1;
  reg L2_5_L1a_3_slc_3_itm;
  reg L2_5_L1a_4_slc_3_itm;
  reg pixel_processing_pixel_processing_if_1_nor_itm;
  reg [2:0] pixel_processing_asn_itm;
  reg [31:0] pixel_processing_if_2_asn_itm;
  reg and_12_itm;
  reg asn_itm_1;
  reg else_io_read_in_data_vld_rsc_svs_st_2;
  reg system_input_output_vld_sva_dfm_st_2;
  reg pixel_processing_pixel_processing_if_1_nor_itm_2;
  reg main_stage_0_2;
  reg and_cse;
  wire and_159_cse;
  wire and_163_cse;
  wire and_171_cse;
  wire and_186_cse;
  wire and_192_cse;
  wire and_193_cse;
  wire and_199_cse;
  wire and_190_cse;
  wire and_184_cse;
  wire clip_window_clip_window_and_1_cse_sva;
  wire pixel_processing_if_2_land_lpi_1_dfm;
  wire system_input_land_1_lpi_1_dfm;
  wire system_input_output_vld_sva_dfm_mx1w0;
  wire [2:0] median_max_8_lpi_1_dfm_mx0;
  wire [2:0] median_max2_9_lpi_1_dfm_1_mx0;
  wire [2:0] median_max2_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_0_lpi_1_dfm_1_mx0;
  wire [2:0] median_max_1_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_4_lpi_1_dfm_mx0;
  wire [2:0] median_max2_8_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_3_lpi_1_dfm_mx0;
  wire [2:0] median_max2_5_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_9_lpi_1_dfm_mx0;
  wire [2:0] median_max2_4_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_6_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_7_1_lpi_1_dfm_mx0;
  wire [2:0] median_max_5_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_6_1_lpi_1_dfm_mx0;
  wire [2:0] pixel_processing_window_6_lpi_1_dfm_mx0;
  wire [2:0] buffer_qr_1_lpi_1_dfm_mx0;
  wire [2:0] buffer_qr_lpi_1_dfm_mx0;
  wire [2:0] median_max2_0_lpi_1_dfm_mx0;
  wire [2:0] median_max_3_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_1_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_4_1_lpi_1_dfm_mx0;
  wire [2:0] clip_window_qr_lpi_1_dfm_mx0;
  wire [2:0] pixel_processing_window_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_6_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_7_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_7_1_lpi_1_dfm_mx0;
  wire [2:0] median_max_8_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_8_1_lpi_1_dfm_mx0;
  wire [2:0] pixel_processing_window_8_lpi_1_dfm_mx0;
  wire [2:0] clip_window_qr_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_1_1_lpi_1_dfm_mx0;
  wire [2:0] median_max_2_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_2_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_3_1_lpi_1_dfm_mx0;
  wire [2:0] pixel_processing_window_0_lpi_1_dfm_mx0;
  wire [2:0] clip_window_qr_3_lpi_1_dfm_mx0;
  wire reg_system_input_system_input_output_vld_and_cse;
  wire and_146_cse;
  wire or_62_cse;
  wire mcu_data_rsci_adr_d_mx0c2;
  wire mcu_data_rsci_adr_d_mx0c3;
  wire [2:0] median_max_5_lpi_1_dfm_mx0;
  wire L1a_if_slc_L1a_if_acc_12_3_itm;
  wire L1b_if_slc_L1b_if_acc_8_3_itm;
  wire L1a_if_slc_L1a_if_acc_9_3_itm;
  wire L1a_if_slc_L1a_if_acc_10_3_itm;
  wire L1b_if_slc_L1b_if_acc_6_3_itm;
  wire L1b_if_slc_L1b_if_acc_3_3_itm;
  wire L1a_if_slc_L1a_if_acc_3_3_itm;
  wire [2:0] L1b_asn_5_mx1w1;
  wire [2:0] L1b_asn_44_mx0w1;
  wire buffer_sel_1_sva_dfm_mx0;
  wire [2:0] median_max2_2_2_lpi_1_dfm_mx0;
  wire [2:0] pixel_processing_mod10_conc_imod_3_1_sva;
  wire [3:0] nl_pixel_processing_mod10_conc_imod_3_1_sva;
  wire [3:0] pixel_processing_mod10_acc_4_psp_sva;
  wire [4:0] nl_pixel_processing_mod10_acc_4_psp_sva;
  wire [5:0] pixel_processing_mod10_acc_psp_sva;
  wire [6:0] nl_pixel_processing_mod10_acc_psp_sva;
  wire [2:0] median_max2_8_lpi_1_dfm_mx0;
  wire [2:0] L1a_asn_13_mx0w1;
  wire [2:0] median_max2_7_lpi_1_dfm_mx0;
  wire [2:0] median_max2_6_3_lpi_1_dfm_mx0;
  wire [2:0] L1a_asn_18_mx0w1;
  wire [2:0] median_max_2_lpi_1_dfm_mx0;
  wire [2:0] median_max2_4_lpi_1_dfm_mx0;
  wire [2:0] median_max_7_2_lpi_1_dfm_mx0;
  wire [2:0] median_max_5_1_lpi_1_dfm_mx0;
  wire [2:0] median_max2_6_lpi_1_dfm_mx0;
  wire [2:0] median_max2_5_lpi_1_dfm_mx0;
  wire L1b_if_acc_11_itm_3;
  wire L1b_if_acc_10_itm_3;
  wire and_133_rgt;
  wire median_max_and_7_rgt;
  wire and_137_rgt;
  wire pixel_processing_and_cse;
  wire reg_median_median_max_or_2_cse;
  wire reg_pixel_processing_pixel_processing_if_1_pixel_processing_if_1_and_cse;
  wire z_out_3;
  wire z_out_1_3;
  wire z_out_2_3;
  wire z_out_3_3;
  wire z_out_4_3;
  wire z_out_5_3;
  wire z_out_6_3;
  wire z_out_7_3;
  wire z_out_8_3;

  wire[7:0] system_input_if_2_qelse_acc_nl;
  wire[8:0] nl_system_input_if_2_qelse_acc_nl;
  wire[0:0] system_input_if_2_system_input_if_2_nand_nl;
  wire[7:0] system_input_if_1_qelse_acc_nl;
  wire[8:0] nl_system_input_if_1_qelse_acc_nl;
  wire[0:0] clip_window_not_6_nl;
  wire[8:0] system_input_else_2_acc_nl;
  wire[9:0] nl_system_input_else_2_acc_nl;
  wire[0:0] system_input_system_input_nand_nl;
  wire[0:0] and_131_nl;
  wire[3:0] L1a_if_acc_15_nl;
  wire[5:0] nl_L1a_if_acc_15_nl;
  wire[2:0] L1b_mux_2_nl;
  wire[2:0] L1b_mux_3_nl;
  wire[0:0] median_max2_and_5_nl;
  wire[0:0] median_max_and_3_nl;
  wire[0:0] median_max2_and_3_nl;
  wire[0:0] median_max_and_1_nl;
  wire[0:0] median_max2_median_max2_nor_nl;
  wire[0:0] buffer_nor_nl;
  wire[0:0] and_147_nl;
  wire[0:0] clip_window_nor_1_nl;
  wire[1:0] pixel_processing_mod10_acc_20_nl;
  wire[2:0] nl_pixel_processing_mod10_acc_20_nl;
  wire[3:0] pixel_processing_mod10_acc_19_nl;
  wire[5:0] nl_pixel_processing_mod10_acc_19_nl;
  wire[5:0] pixel_processing_mod10_acc_18_nl;
  wire[6:0] nl_pixel_processing_mod10_acc_18_nl;
  wire[4:0] pixel_processing_mod10_acc_17_nl;
  wire[5:0] nl_pixel_processing_mod10_acc_17_nl;
  wire[3:0] pixel_processing_mod10_acc_15_nl;
  wire[4:0] nl_pixel_processing_mod10_acc_15_nl;
  wire[2:0] pixel_processing_mod10_acc_11_nl;
  wire[3:0] nl_pixel_processing_mod10_acc_11_nl;
  wire[2:0] pixel_processing_mod10_acc_10_nl;
  wire[3:0] nl_pixel_processing_mod10_acc_10_nl;
  wire[3:0] pixel_processing_mod10_acc_14_nl;
  wire[4:0] nl_pixel_processing_mod10_acc_14_nl;
  wire[2:0] pixel_processing_mod10_acc_9_nl;
  wire[3:0] nl_pixel_processing_mod10_acc_9_nl;
  wire[2:0] pixel_processing_mod10_acc_8_nl;
  wire[3:0] nl_pixel_processing_mod10_acc_8_nl;
  wire[4:0] pixel_processing_mod10_acc_16_nl;
  wire[5:0] nl_pixel_processing_mod10_acc_16_nl;
  wire[3:0] pixel_processing_mod10_acc_13_nl;
  wire[4:0] nl_pixel_processing_mod10_acc_13_nl;
  wire[2:0] pixel_processing_mod10_acc_7_nl;
  wire[3:0] nl_pixel_processing_mod10_acc_7_nl;
  wire[2:0] pixel_processing_mod10_acc_6_nl;
  wire[3:0] nl_pixel_processing_mod10_acc_6_nl;
  wire[3:0] pixel_processing_mod10_acc_12_nl;
  wire[4:0] nl_pixel_processing_mod10_acc_12_nl;
  wire[2:0] pixel_processing_mod10_acc_5_nl;
  wire[3:0] nl_pixel_processing_mod10_acc_5_nl;
  wire[3:0] L1b_if_acc_7_nl;
  wire[5:0] nl_L1b_if_acc_7_nl;
  wire[3:0] L1b_if_acc_11_nl;
  wire[5:0] nl_L1b_if_acc_11_nl;
  wire[3:0] L1b_if_acc_10_nl;
  wire[5:0] nl_L1b_if_acc_10_nl;
  wire[0:0] nand_nl;
  wire[3:0] L1a_if_acc_12_nl;
  wire[5:0] nl_L1a_if_acc_12_nl;
  wire[3:0] L1b_if_acc_8_nl;
  wire[5:0] nl_L1b_if_acc_8_nl;
  wire[3:0] L1a_if_acc_9_nl;
  wire[5:0] nl_L1a_if_acc_9_nl;
  wire[3:0] L1a_if_acc_10_nl;
  wire[5:0] nl_L1a_if_acc_10_nl;
  wire[3:0] L1b_if_acc_6_nl;
  wire[5:0] nl_L1b_if_acc_6_nl;
  wire[3:0] L1b_if_acc_3_nl;
  wire[5:0] nl_L1b_if_acc_3_nl;
  wire[3:0] L1a_if_acc_3_nl;
  wire[5:0] nl_L1a_if_acc_3_nl;
  wire[0:0] system_input_c_system_input_c_or_nl;
  wire[2:0] system_input_c_and_nl;
  wire[2:0] system_input_c_mux1h_nl;
  wire[0:0] system_input_c_nor_1_nl;
  wire[31:0] pixel_processing_if_2_mux1h_nl;
  wire[31:0] pixel_processing_if_1_pixel_processing_if_1_acc_1_nl;
  wire[32:0] nl_pixel_processing_if_1_pixel_processing_if_1_acc_1_nl;
  wire[0:0] or_149_nl;
  wire[0:0] mcu_data_nor_nl;
  wire[9:0] buffer_buf_mux_3_nl;
  wire[0:0] buffer_buf_nor_nl;
  wire[9:0] buffer_buf_mux_2_nl;
  wire[0:0] buffer_buf_nor_1_nl;
  wire[4:0] acc_nl;
  wire[5:0] nl_acc_nl;
  wire[2:0] thresholding_if_mux1h_3_nl;
  wire[0:0] thresholding_if_and_2_nl;
  wire[0:0] thresholding_if_and_3_nl;
  wire[2:0] thresholding_if_mux1h_4_nl;
  wire[2:0] L1b_mux_30_nl;
  wire[4:0] acc_1_nl;
  wire[5:0] nl_acc_1_nl;
  wire[2:0] L1a_if_mux_19_nl;
  wire[2:0] L1a_if_mux_20_nl;
  wire[4:0] acc_2_nl;
  wire[5:0] nl_acc_2_nl;
  wire[2:0] L1a_if_mux_21_nl;
  wire[2:0] L1a_if_mux_22_nl;
  wire[4:0] acc_3_nl;
  wire[5:0] nl_acc_3_nl;
  wire[2:0] L1b_if_mux1h_3_nl;
  wire[2:0] L1b_if_mux1h_4_nl;
  wire[4:0] acc_4_nl;
  wire[5:0] nl_acc_4_nl;
  wire[2:0] L1b_if_mux_6_nl;
  wire[2:0] L1b_if_mux_7_nl;
  wire[4:0] acc_5_nl;
  wire[5:0] nl_acc_5_nl;
  wire[2:0] L1a_if_mux_23_nl;
  wire[2:0] L1a_if_mux_24_nl;
  wire[2:0] clip_window_mux_8_nl;
  wire[4:0] acc_6_nl;
  wire[5:0] nl_acc_6_nl;
  wire[2:0] L1a_if_mux_25_nl;
  wire[2:0] L1a_if_mux_26_nl;
  wire[4:0] acc_7_nl;
  wire[5:0] nl_acc_7_nl;
  wire[2:0] L1b_if_mux_8_nl;
  wire[2:0] L1b_if_mux_9_nl;
  wire[4:0] acc_8_nl;
  wire[5:0] nl_acc_8_nl;
  wire[2:0] L1a_if_mux_27_nl;
  wire[2:0] L1a_if_mux_28_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [2:0] nl_out_data_rsci_d;
  assign nl_out_data_rsci_d = {{2{out_data_rsci_d_0}}, out_data_rsci_d_0};
  wire [0:0] nl_filter_core_core_fsm_inst_buffer_buf_vinit_C_1_tr0;
  assign nl_filter_core_core_fsm_inst_buffer_buf_vinit_C_1_tr0 = ~ buffer_buf_buffer_buf_nor_itm_1;
  mgc_in_wire_en_v1 #(.rscid(32'sd1),
  .width(32'sd3)) in_data_rsci (
      .ld(in_data_rsci_ld),
      .d(in_data_rsci_d),
      .lz(in_data_rsc_lz),
      .z(in_data_rsc_z)
    );
  mgc_in_wire_v1 #(.rscid(32'sd2),
  .width(32'sd1)) in_data_vld_rsci (
      .d(in_data_vld_rsci_d),
      .z(in_data_vld_rsc_z)
    );
  mgc_out_stdreg_en_v1 #(.rscid(32'sd3),
  .width(32'sd3)) out_data_rsci (
      .ld(out_data_rsci_ld),
      .d(nl_out_data_rsci_d[2:0]),
      .lz(out_data_rsc_lz),
      .z(out_data_rsc_z)
    );
  filter_core_core_fsm filter_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .buffer_buf_vinit_C_1_tr0(nl_filter_core_core_fsm_inst_buffer_buf_vinit_C_1_tr0[0:0])
    );
  assign or_62_cse = or_dcpl_1 | (~ (fsm_output[3]));
  assign reg_system_input_system_input_output_vld_and_cse = in_data_vld_rsci_d &
      mcu_ready_sva & (fsm_output[3]);
  assign reg_pixel_processing_pixel_processing_if_1_pixel_processing_if_1_and_cse
      = mcu_ready_sva & (~ or_tmp_49);
  assign pixel_processing_and_cse = mcu_ready_sva & (fsm_output[5]);
  assign and_133_rgt = mcu_ready_sva & (~ z_out_3_3) & (fsm_output[5]);
  assign median_max_and_7_rgt = mcu_ready_sva & (~ L1b_if_acc_11_itm_3) & (fsm_output[5]);
  assign reg_median_median_max_or_2_cse = (mcu_ready_sva & L1b_if_acc_11_itm_3 &
      (fsm_output[5])) | median_max_and_7_rgt;
  assign and_137_rgt = mcu_ready_sva & (~ L1b_if_acc_10_itm_3) & (fsm_output[5]);
  assign and_146_cse = (system_input_r_filter_sva==8'b11101111);
  assign L1b_asn_5_mx1w1 = MUX_v_3_2_2(L1a_asn_18_mx0w1, median_max_5_1_lpi_1_dfm_mx0,
      L1a_if_slc_L1a_if_acc_12_3_itm);
  assign median_max_5_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_6_lpi_1_dfm_mx0, median_max2_5_lpi_1_dfm_mx0,
      z_out_3_3);
  assign system_input_output_vld_sva_dfm_mx1w0 = system_input_output_vld_sva | ((system_input_c_sva==9'b000000001)
      & (system_input_r_sva==8'b00000001));
  assign pixel_processing_if_2_land_lpi_1_dfm = ((pixel_processing_frame_sva[31:1]!=31'b0000000000000000000000000000000))
      & (pixel_processing_frame_sva[0]) & (pixel_processing_mod10_acc_3_tmp==3'b000);
  assign system_input_land_1_lpi_1_dfm = clip_window_clip_window_and_1_cse_sva &
      and_146_cse;
  assign L1b_asn_44_mx0w1 = MUX_v_3_2_2(median_max2_0_lpi_1_dfm_mx0, median_max_1_1_lpi_1_dfm_mx0,
      z_out_6_3);
  assign clip_window_clip_window_and_1_cse_sva = (system_input_c_filter_sva==9'b100111111);
  assign buffer_nor_nl = ~((system_input_c_sva!=9'b000000000));
  assign buffer_sel_1_sva_dfm_mx0 = MUX_s_1_2_2(buffer_sel_1_sva, (~ buffer_sel_1_sva),
      buffer_nor_nl);
  assign nl_pixel_processing_mod10_acc_3_tmp = conv_u2u_1_3(pixel_processing_mod10_conc_imod_3_1_sva[2])
      + conv_u2u_2_3(pixel_processing_mod10_conc_imod_3_1_sva[1:0]);
  assign pixel_processing_mod10_acc_3_tmp = nl_pixel_processing_mod10_acc_3_tmp[2:0];
  assign median_max2_0_lpi_1_dfm_1_mx0 = MUX_v_3_2_2(median_max_1_1_lpi_1_dfm_mx0,
      median_max2_0_lpi_1_dfm_mx0, z_out_6_3);
  assign median_max_1_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_2_2_lpi_1_dfm_mx0,
      L1b_asn_44_mx0w1, z_out_3_3);
  assign median_max2_2_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_3_1_lpi_1_dfm_mx0,
      median_max_2_1_lpi_1_dfm_mx0, z_out_2_3);
  assign median_max_2_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_1_1_lpi_1_dfm_mx0,
      median_max2_2_1_lpi_1_dfm_mx0, z_out_7_3);
  assign median_max_3_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_4_1_lpi_1_dfm_mx0,
      median_max2_3_1_lpi_1_dfm_mx0, z_out_4_3);
  assign median_max2_0_lpi_1_dfm_mx0 = MUX_v_3_2_2(clip_window_qr_lpi_1_dfm_mx0,
      pixel_processing_window_0_lpi_1_dfm_mx0, z_out_8_3);
  assign median_max_1_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_2_1_lpi_1_dfm_mx0,
      median_max2_1_1_lpi_1_dfm_mx0, z_out_7_3);
  assign median_max2_3_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(pixel_processing_window_2_lpi_1_dfm_mx0,
      clip_window_qr_3_lpi_1_dfm_mx0, z_out_1_3);
  assign and_147_nl = or_dcpl_124 & (~ z_out_5_3);
  assign median_max2_4_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_window_7_sva, system_input_window_8_sva,
      and_147_nl);
  assign median_max2_1_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(pixel_processing_window_0_lpi_1_dfm_mx0,
      clip_window_qr_lpi_1_dfm_mx0, z_out_8_3);
  assign median_max2_2_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(clip_window_qr_3_lpi_1_dfm_mx0,
      pixel_processing_window_2_lpi_1_dfm_mx0, z_out_1_3);
  assign pixel_processing_window_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_window_4_sva,
      system_input_window_5_sva, or_dcpl_124);
  assign clip_window_qr_3_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_window_6_sva,
      system_input_window_7_sva, and_dcpl_126);
  assign pixel_processing_window_0_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_window_3_sva,
      system_input_window_4_sva, and_dcpl_126);
  assign clip_window_nor_1_nl = ~((system_input_c_filter_sva!=9'b000000000));
  assign clip_window_qr_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_window_4_sva, system_input_window_7_sva,
      clip_window_nor_1_nl);
  assign nl_pixel_processing_mod10_acc_20_nl = conv_s2s_1_2(~ (pixel_processing_mod10_acc_4_psp_sva[3]))
      + conv_u2s_1_2(~ (pixel_processing_mod10_acc_4_psp_sva[2]));
  assign pixel_processing_mod10_acc_20_nl = nl_pixel_processing_mod10_acc_20_nl[1:0];
  assign nl_pixel_processing_mod10_conc_imod_3_1_sva = conv_s2u_2_3(pixel_processing_mod10_acc_20_nl)
      + ({(pixel_processing_mod10_acc_4_psp_sva[3]) , (pixel_processing_mod10_acc_4_psp_sva[1:0])});
  assign pixel_processing_mod10_conc_imod_3_1_sva = nl_pixel_processing_mod10_conc_imod_3_1_sva[2:0];
  assign nl_pixel_processing_mod10_acc_19_nl = conv_u2s_2_4(~ (pixel_processing_mod10_acc_psp_sva[3:2]))
      + conv_s2s_2_4(pixel_processing_mod10_acc_psp_sva[5:4]) + 4'b1;
  assign pixel_processing_mod10_acc_19_nl = nl_pixel_processing_mod10_acc_19_nl[3:0];
  assign nl_pixel_processing_mod10_acc_4_psp_sva = (pixel_processing_mod10_acc_19_nl)
      + conv_s2u_3_4({1'b1 , (pixel_processing_mod10_acc_psp_sva[1:0])});
  assign pixel_processing_mod10_acc_4_psp_sva = nl_pixel_processing_mod10_acc_4_psp_sva[3:0];
  assign nl_pixel_processing_mod10_acc_11_nl = conv_u2u_2_3(~ (pixel_processing_frame_sva[4:3]))
      + conv_u2u_2_3(pixel_processing_frame_sva[6:5]);
  assign pixel_processing_mod10_acc_11_nl = nl_pixel_processing_mod10_acc_11_nl[2:0];
  assign nl_pixel_processing_mod10_acc_10_nl = conv_u2u_2_3(~ (pixel_processing_frame_sva[8:7]))
      + conv_u2u_2_3(pixel_processing_frame_sva[10:9]);
  assign pixel_processing_mod10_acc_10_nl = nl_pixel_processing_mod10_acc_10_nl[2:0];
  assign nl_pixel_processing_mod10_acc_15_nl = conv_u2u_3_4(pixel_processing_mod10_acc_11_nl)
      + conv_u2u_3_4(pixel_processing_mod10_acc_10_nl);
  assign pixel_processing_mod10_acc_15_nl = nl_pixel_processing_mod10_acc_15_nl[3:0];
  assign nl_pixel_processing_mod10_acc_9_nl = conv_u2u_2_3(~ (pixel_processing_frame_sva[12:11]))
      + conv_u2u_2_3(pixel_processing_frame_sva[14:13]);
  assign pixel_processing_mod10_acc_9_nl = nl_pixel_processing_mod10_acc_9_nl[2:0];
  assign nl_pixel_processing_mod10_acc_8_nl = conv_u2u_2_3(~ (pixel_processing_frame_sva[16:15]))
      + conv_u2u_2_3(pixel_processing_frame_sva[18:17]);
  assign pixel_processing_mod10_acc_8_nl = nl_pixel_processing_mod10_acc_8_nl[2:0];
  assign nl_pixel_processing_mod10_acc_14_nl = conv_u2u_3_4(pixel_processing_mod10_acc_9_nl)
      + conv_u2u_3_4(pixel_processing_mod10_acc_8_nl);
  assign pixel_processing_mod10_acc_14_nl = nl_pixel_processing_mod10_acc_14_nl[3:0];
  assign nl_pixel_processing_mod10_acc_17_nl = conv_u2u_4_5(pixel_processing_mod10_acc_15_nl)
      + conv_u2u_4_5(pixel_processing_mod10_acc_14_nl);
  assign pixel_processing_mod10_acc_17_nl = nl_pixel_processing_mod10_acc_17_nl[4:0];
  assign nl_pixel_processing_mod10_acc_7_nl = conv_u2u_2_3(~ (pixel_processing_frame_sva[20:19]))
      + conv_u2u_2_3(pixel_processing_frame_sva[22:21]);
  assign pixel_processing_mod10_acc_7_nl = nl_pixel_processing_mod10_acc_7_nl[2:0];
  assign nl_pixel_processing_mod10_acc_6_nl = conv_u2u_2_3(~ (pixel_processing_frame_sva[24:23]))
      + conv_u2u_2_3(pixel_processing_frame_sva[26:25]);
  assign pixel_processing_mod10_acc_6_nl = nl_pixel_processing_mod10_acc_6_nl[2:0];
  assign nl_pixel_processing_mod10_acc_13_nl = conv_u2u_3_4(pixel_processing_mod10_acc_7_nl)
      + conv_u2u_3_4(pixel_processing_mod10_acc_6_nl);
  assign pixel_processing_mod10_acc_13_nl = nl_pixel_processing_mod10_acc_13_nl[3:0];
  assign nl_pixel_processing_mod10_acc_5_nl = conv_u2u_2_3(~ (pixel_processing_frame_sva[28:27]))
      + conv_u2u_2_3(pixel_processing_frame_sva[30:29]);
  assign pixel_processing_mod10_acc_5_nl = nl_pixel_processing_mod10_acc_5_nl[2:0];
  assign nl_pixel_processing_mod10_acc_12_nl = conv_u2u_3_4(pixel_processing_mod10_acc_5_nl)
      + conv_u2u_2_4(pixel_processing_frame_sva[2:1]);
  assign pixel_processing_mod10_acc_12_nl = nl_pixel_processing_mod10_acc_12_nl[3:0];
  assign nl_pixel_processing_mod10_acc_16_nl = conv_u2u_4_5(pixel_processing_mod10_acc_13_nl)
      + conv_u2u_4_5(pixel_processing_mod10_acc_12_nl);
  assign pixel_processing_mod10_acc_16_nl = nl_pixel_processing_mod10_acc_16_nl[4:0];
  assign nl_pixel_processing_mod10_acc_18_nl = conv_u2u_5_6(pixel_processing_mod10_acc_17_nl)
      + conv_u2u_5_6(pixel_processing_mod10_acc_16_nl);
  assign pixel_processing_mod10_acc_18_nl = nl_pixel_processing_mod10_acc_18_nl[5:0];
  assign nl_pixel_processing_mod10_acc_psp_sva = (pixel_processing_mod10_acc_18_nl)
      + ({5'b10101 , (~ (pixel_processing_frame_sva[31]))});
  assign pixel_processing_mod10_acc_psp_sva = nl_pixel_processing_mod10_acc_psp_sva[5:0];
  assign and_tmp = in_data_vld_rsci_d & mcu_ready_sva;
  assign if_if_if_and_tmp = (mcu_data_rsci_q_d==32'b00000000000000000000000000000001);
  assign median_max2_8_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_9_lpi_1_dfm_1_mx0,
      median_max_8_lpi_1_dfm_mx0, z_out_2_3);
  assign L1a_asn_13_mx0w1 = MUX_v_3_2_2(median_max_4_lpi_1_dfm_mx0, median_max2_6_2_lpi_1_dfm_mx0,
      L1b_if_slc_L1b_if_acc_8_3_itm);
  assign median_max2_7_lpi_1_dfm_mx0 = MUX_v_3_2_2(L1a_asn_13_mx0w1, median_max_7_2_lpi_1_dfm_mx0,
      z_out_6_3);
  assign median_max2_6_3_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_7_2_lpi_1_dfm_mx0,
      L1a_asn_13_mx0w1, z_out_6_3);
  assign L1a_asn_18_mx0w1 = MUX_v_3_2_2(median_max_2_2_lpi_1_dfm, median_max_3_lpi_1_dfm_mx0,
      L1a_if_slc_L1a_if_acc_9_3_itm);
  assign nl_L1b_if_acc_7_nl = ({1'b1 , median_max2_1_lpi_1_dfm}) + conv_u2u_3_4(~
      median_max2_2_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_7_nl = nl_L1b_if_acc_7_nl[3:0];
  assign median_max_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_1_lpi_1_dfm, median_max2_2_lpi_1_dfm_mx0,
      readslicef_4_1_3((L1b_if_acc_7_nl)));
  assign median_max2_4_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_5_1_lpi_1_dfm_mx0,
      L1a_asn_18_mx0w1, L1a_if_slc_L1a_if_acc_12_3_itm);
  assign median_max2_9_lpi_1_dfm_1_mx0 = MUX_v_3_2_2(median_max_8_1_lpi_1_dfm_mx0,
      median_max2_9_lpi_1_dfm_mx0, z_out_8_3);
  assign median_max_8_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_7_2_lpi_1_dfm_mx0,
      median_max2_8_2_lpi_1_dfm_mx0, z_out_7_3);
  assign median_max_7_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_8_2_lpi_1_dfm_mx0,
      median_max2_7_2_lpi_1_dfm_mx0, z_out_7_3);
  assign median_max_5_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_6_2_lpi_1_dfm_mx0,
      median_max_4_lpi_1_dfm_mx0, L1b_if_slc_L1b_if_acc_8_3_itm);
  assign median_max2_8_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_9_lpi_1_dfm_mx0,
      median_max_8_1_lpi_1_dfm_mx0, z_out_8_3);
  assign median_max2_7_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_5_2_lpi_1_dfm_mx0,
      median_max_7_1_lpi_1_dfm_mx0, L1a_if_slc_L1a_if_acc_10_3_itm);
  assign median_max_4_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_3_2_lpi_1_dfm, median_max2_4_2_lpi_1_dfm_mx0,
      z_out_4_3);
  assign median_max2_6_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_7_1_lpi_1_dfm_mx0,
      median_max2_5_2_lpi_1_dfm_mx0, L1a_if_slc_L1a_if_acc_10_3_itm);
  assign median_max2_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_3_lpi_1_dfm_mx0, median_max_2_2_lpi_1_dfm,
      L1a_if_slc_L1a_if_acc_9_3_itm);
  assign median_max2_9_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_7_1_lpi_1_dfm_mx0,
      pixel_processing_window_8_lpi_1_dfm_mx0, z_out_5_3);
  assign median_max_8_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_6_2_lpi_1_dfm_mx0,
      median_max2_8_1_lpi_1_dfm_mx0, L1b_if_slc_L1b_if_acc_6_3_itm);
  assign median_max2_5_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_4_2_lpi_1_dfm, median_max_5_2_lpi_1_dfm_mx0,
      z_out_1_3);
  assign median_max_7_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_8_1_lpi_1_dfm_mx0,
      median_max_6_2_lpi_1_dfm_mx0, L1b_if_slc_L1b_if_acc_6_3_itm);
  assign median_max_3_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_4_2_lpi_1_dfm_mx0,
      median_max2_3_2_lpi_1_dfm, z_out_4_3);
  assign median_max_6_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_5_1_lpi_1_dfm, median_max2_6_1_lpi_1_dfm_mx0,
      L1b_if_slc_L1b_if_acc_3_3_itm);
  assign median_max2_8_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(pixel_processing_window_8_lpi_1_dfm_mx0,
      median_max2_7_1_lpi_1_dfm_mx0, z_out_5_3);
  assign median_max2_4_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_5_2_lpi_1_dfm_mx0,
      median_max_4_2_lpi_1_dfm, z_out_1_3);
  assign pixel_processing_window_8_lpi_1_dfm_mx0 = MUX_v_3_2_2(system_input_din_sva_1,
      buffer_qr_1_lpi_1_dfm_mx0, clip_window_ac_int_cctor_2_sva_1);
  assign median_max2_7_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(pixel_processing_window_6_lpi_1_dfm_mx0,
      clip_window_qr_2_lpi_1_dfm_mx0, L1a_if_slc_L1a_if_acc_3_3_itm);
  assign median_max_5_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max2_6_1_lpi_1_dfm_mx0,
      median_max2_5_1_lpi_1_dfm, L1b_if_slc_L1b_if_acc_3_3_itm);
  assign median_max2_6_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(clip_window_qr_2_lpi_1_dfm_mx0,
      pixel_processing_window_6_lpi_1_dfm_mx0, L1a_if_slc_L1a_if_acc_3_3_itm);
  assign pixel_processing_window_6_lpi_1_dfm_mx0 = MUX_v_3_2_2(buffer_qr_1_lpi_1_dfm_mx0,
      buffer_qr_lpi_1_dfm_mx0, clip_window_unequal_tmp_2);
  assign clip_window_qr_2_lpi_1_dfm_mx0 = MUX_v_3_2_2(buffer_qr_1_lpi_1_dfm_mx0,
      system_input_window_7_sva, clip_window_clip_window_and_1_cse_sva_1);
  assign buffer_qr_1_lpi_1_dfm_mx0 = MUX_v_3_2_2(buffer_buf_rsci_q_d, buffer_t0_sva_1,
      buffer_sel_1_sva_dfm);
  assign buffer_qr_lpi_1_dfm_mx0 = MUX_v_3_2_2(buffer_t0_sva_1, buffer_buf_rsci_q_d,
      buffer_sel_1_sva_dfm);
  assign median_max2_6_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_7_lpi_1_dfm, median_max_6_lpi_1_dfm,
      L2_5_L1a_4_slc_3_itm);
  assign median_max2_5_lpi_1_dfm_mx0 = MUX_v_3_2_2(median_max_4_1_lpi_1_dfm, median_max_5_3_lpi_1_dfm,
      L2_5_L1a_3_slc_3_itm);
  assign nl_L1b_if_acc_11_nl = ({1'b1 , L1b_asn_5_mx1w1}) + conv_u2u_3_4(~ median_max2_6_3_lpi_1_dfm_mx0)
      + 4'b1;
  assign L1b_if_acc_11_nl = nl_L1b_if_acc_11_nl[3:0];
  assign L1b_if_acc_11_itm_3 = readslicef_4_1_3((L1b_if_acc_11_nl));
  assign nl_L1b_if_acc_10_nl = ({1'b1 , median_max_2_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max2_4_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_10_nl = nl_L1b_if_acc_10_nl[3:0];
  assign L1b_if_acc_10_itm_3 = readslicef_4_1_3((L1b_if_acc_10_nl));
  assign or_dcpl_1 = ~(in_data_vld_rsci_d & mcu_ready_sva);
  assign and_dcpl_41 = else_io_read_in_data_vld_rsc_svs & system_input_output_vld_sva_dfm;
  assign or_dcpl_54 = ~(else_io_read_in_data_vld_rsc_svs & system_input_output_vld_sva_dfm);
  assign nor_tmp_5 = system_input_land_1_lpi_1_dfm_1 & system_input_output_vld_sva_dfm
      & else_io_read_in_data_vld_rsc_svs;
  assign nor_tmp_6 = mcu_ready_sva & system_input_land_1_lpi_1_dfm_1 & system_input_output_vld_sva_dfm
      & else_io_read_in_data_vld_rsc_svs;
  assign nand_nl = ~(mcu_ready_sva & (~ nor_tmp_5));
  assign mux_tmp_6 = MUX_s_1_2_2(nor_tmp_6, (nand_nl), if_if_if_and_tmp);
  assign or_dcpl_75 = (system_input_c_sva[7]) | (system_input_c_sva[6]) | (~ (system_input_c_sva[0]));
  assign or_dcpl_80 = ~((system_input_r_filter_sva[3]) & (system_input_r_filter_sva[5])
      & (system_input_r_filter_sva[6]) & (system_input_r_filter_sva[7]));
  assign or_dcpl_81 = ~((system_input_r_filter_sva[2:1]==2'b11));
  assign or_dcpl_87 = ~((system_input_c_filter_sva[5:4]==2'b11));
  assign and_dcpl_101 = ~((~(or_dcpl_75 | (system_input_c_sva[8]) | (system_input_c_sva[5])
      | (system_input_c_sva[4]) | (system_input_c_sva[3]) | (system_input_c_sva[2])
      | (system_input_c_sva[1]) | (system_input_r_sva!=8'b00000001))) | system_input_output_vld_sva);
  assign or_dcpl_124 = (system_input_r_filter_sva[4]) | (~ (system_input_r_filter_sva[0]))
      | or_dcpl_81 | or_dcpl_80;
  assign and_dcpl_126 = ~((system_input_r_filter_sva!=8'b00000000));
  assign nl_L1a_if_acc_12_nl = ({1'b1 , L1a_asn_18_mx0w1}) + conv_u2u_3_4(~ median_max_5_1_lpi_1_dfm_mx0)
      + 4'b1;
  assign L1a_if_acc_12_nl = nl_L1a_if_acc_12_nl[3:0];
  assign L1a_if_slc_L1a_if_acc_12_3_itm = readslicef_4_1_3((L1a_if_acc_12_nl));
  assign nl_L1b_if_acc_8_nl = ({1'b1 , median_max_4_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max2_6_2_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_8_nl = nl_L1b_if_acc_8_nl[3:0];
  assign L1b_if_slc_L1b_if_acc_8_3_itm = readslicef_4_1_3((L1b_if_acc_8_nl));
  assign nl_L1a_if_acc_9_nl = ({1'b1 , median_max_2_2_lpi_1_dfm}) + conv_u2u_3_4(~
      median_max_3_lpi_1_dfm_mx0) + 4'b1;
  assign L1a_if_acc_9_nl = nl_L1a_if_acc_9_nl[3:0];
  assign L1a_if_slc_L1a_if_acc_9_3_itm = readslicef_4_1_3((L1a_if_acc_9_nl));
  assign nl_L1a_if_acc_10_nl = ({1'b1 , median_max2_5_2_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max_7_1_lpi_1_dfm_mx0) + 4'b1;
  assign L1a_if_acc_10_nl = nl_L1a_if_acc_10_nl[3:0];
  assign L1a_if_slc_L1a_if_acc_10_3_itm = readslicef_4_1_3((L1a_if_acc_10_nl));
  assign nl_L1b_if_acc_6_nl = ({1'b1 , median_max_6_2_lpi_1_dfm_mx0}) + conv_u2u_3_4(~
      median_max2_8_1_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_6_nl = nl_L1b_if_acc_6_nl[3:0];
  assign L1b_if_slc_L1b_if_acc_6_3_itm = readslicef_4_1_3((L1b_if_acc_6_nl));
  assign nl_L1b_if_acc_3_nl = ({1'b1 , median_max2_5_1_lpi_1_dfm}) + conv_u2u_3_4(~
      median_max2_6_1_lpi_1_dfm_mx0) + 4'b1;
  assign L1b_if_acc_3_nl = nl_L1b_if_acc_3_nl[3:0];
  assign L1b_if_slc_L1b_if_acc_3_3_itm = readslicef_4_1_3((L1b_if_acc_3_nl));
  assign nl_L1a_if_acc_3_nl = ({1'b1 , pixel_processing_window_6_lpi_1_dfm_mx0})
      + conv_u2u_3_4(~ clip_window_qr_2_lpi_1_dfm_mx0) + 4'b1;
  assign L1a_if_acc_3_nl = nl_L1a_if_acc_3_nl[3:0];
  assign L1a_if_slc_L1a_if_acc_3_3_itm = readslicef_4_1_3((L1a_if_acc_3_nl));
  assign and_159_cse = and_tmp & (fsm_output[3]);
  assign and_163_cse = else_io_read_in_data_vld_rsc_svs & mcu_ready_sva & (fsm_output[4]);
  assign and_171_cse = (~(else_io_read_in_data_vld_rsc_svs & mcu_ready_sva)) & (fsm_output[4]);
  assign and_184_cse = and_dcpl_41 & asn_itm & pixel_processing_pixel_processing_if_1_nor_itm
      & (fsm_output[6]);
  assign and_186_cse = pixel_processing_pixel_processing_if_1_nor_itm_2 & system_input_output_vld_sva_dfm_st_2
      & else_io_read_in_data_vld_rsc_svs_st_2 & asn_itm_1 & main_stage_0_2 & (fsm_output[3]);
  assign and_190_cse = nor_tmp_6 & (fsm_output[5]);
  assign and_192_cse = ((~(pixel_processing_pixel_processing_if_1_nor_itm_2 & system_input_output_vld_sva_dfm_st_2
      & else_io_read_in_data_vld_rsc_svs_st_2)) | (~(asn_itm_1 & main_stage_0_2)))
      & (fsm_output[3]);
  assign and_193_cse = (~ mux_tmp_6) & (fsm_output[5]);
  assign and_199_cse = (~ mcu_ready_sva) & if_if_if_and_tmp & (fsm_output[5]);
  assign or_tmp_35 = and_cse & (fsm_output[5]);
  assign or_tmp_49 = (fsm_output[5:4]!=2'b00);
  assign mcu_data_rsci_adr_d_mx0c2 = and_199_cse | ((~ mcu_ready_sva) & (fsm_output[4]));
  assign mcu_data_rsci_adr_d_mx0c3 = nor_tmp_5 & mcu_ready_sva & pixel_processing_if_2_land_lpi_1_dfm_1
      & (fsm_output[4]);
  assign system_input_c_system_input_c_or_nl = mcu_data_rsci_adr_d_mx0c2 | mcu_data_rsci_adr_d_mx0c3
      | and_190_cse;
  assign system_input_c_mux1h_nl = MUX1HOT_v_3_4_2(median_max_5_lpi_1_dfm_5, 3'b1,
      3'b10, median_max_5_lpi_1_dfm_mx0, {and_186_cse , mcu_data_rsci_adr_d_mx0c3
      , and_190_cse , and_184_cse});
  assign system_input_c_nor_1_nl = ~(and_192_cse | and_193_cse | (fsm_output[2:0]!=3'b000)
      | ((or_dcpl_54 | (~(asn_itm & pixel_processing_pixel_processing_if_1_nor_itm)))
      & (fsm_output[6])) | ((or_dcpl_54 | (~(system_input_land_1_lpi_1_dfm_1 & pixel_processing_if_2_land_lpi_1_dfm_1)))
      & mcu_ready_sva & (fsm_output[4])) | mcu_data_rsci_adr_d_mx0c2);
  assign system_input_c_and_nl = MUX_v_3_2_2(3'b000, (system_input_c_mux1h_nl), (system_input_c_nor_1_nl));
  assign mcu_data_rsci_adr_d = {5'b0 , (system_input_c_system_input_c_or_nl) , (system_input_c_and_nl)};
  assign nl_pixel_processing_if_1_pixel_processing_if_1_acc_1_nl = mcu_data_rsci_q_d
      + 32'b1;
  assign pixel_processing_if_1_pixel_processing_if_1_acc_1_nl = nl_pixel_processing_if_1_pixel_processing_if_1_acc_1_nl[31:0];
  assign or_149_nl = and_190_cse | (fsm_output[0]);
  assign pixel_processing_if_2_mux1h_nl = MUX1HOT_v_32_3_2(pixel_processing_if_2_asn_itm,
      (pixel_processing_if_1_pixel_processing_if_1_acc_1_nl), 32'b10, {(or_149_nl)
      , and_186_cse , and_199_cse});
  assign mcu_data_nor_nl = ~(and_192_cse | and_193_cse | (~((fsm_output[0]) | (fsm_output[5])
      | (fsm_output[3]))));
  assign mcu_data_rsci_d_d = MUX_v_32_2_2(32'b00000000000000000000000000000000, (pixel_processing_if_2_mux1h_nl),
      (mcu_data_nor_nl));
  assign mcu_data_rsci_we_d = and_186_cse | (mux_tmp_6 & (fsm_output[5]));
  assign mcu_data_rsci_ram_rw_A_internal_RMASK_B_d = and_184_cse | ((~((~(and_dcpl_41
      & system_input_land_1_lpi_1_dfm_1 & pixel_processing_if_2_land_lpi_1_dfm_1))
      & mcu_ready_sva)) & (fsm_output[4]));
  assign buffer_buf_mux_3_nl = MUX_v_10_2_2(({1'b0 , system_input_c_sva}), ({buffer_acc_1_itm_2
      , buffer_slc_buffer_c_5_0_1_itm_2}), and_163_cse);
  assign buffer_buf_nor_nl = ~((or_dcpl_1 & (fsm_output[3])) | (~((fsm_output[4:3]!=2'b00)))
      | and_171_cse);
  assign buffer_buf_rsci_radr_d = MUX_v_10_2_2(10'b0000000000, (buffer_buf_mux_3_nl),
      (buffer_buf_nor_nl));
  assign buffer_buf_mux_2_nl = MUX_v_10_2_2(buffer_buf_vinit_ndx_sva, ({buffer_acc_3_itm_2
      , buffer_slc_buffer_c_5_0_1_itm_2}), and_163_cse);
  assign buffer_buf_nor_1_nl = ~((~((fsm_output[1]) | (fsm_output[4]))) | and_171_cse);
  assign buffer_buf_rsci_wadr_d = MUX_v_10_2_2(10'b0000000000, (buffer_buf_mux_2_nl),
      (buffer_buf_nor_1_nl));
  assign buffer_buf_rsci_d_d = MUX_v_3_2_2(3'b000, in_data_rsci_d, and_163_cse);
  assign buffer_buf_rsci_we_d = (fsm_output[1]) | and_163_cse;
  assign buffer_buf_rsci_re_d = and_159_cse | and_163_cse;
  always @(posedge clk) begin
    if ( rst ) begin
      out_data_rsci_d_0 <= 1'b0;
    end
    else if ( ~((~ (fsm_output[6])) | or_dcpl_54 | (~ asn_itm)) ) begin
      out_data_rsci_d_0 <= ~ z_out_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      out_data_rsci_ld <= 1'b0;
      in_data_rsci_ld <= 1'b0;
      buffer_buf_buffer_buf_nor_itm_1 <= 1'b0;
      buffer_buf_acc_itm_2 <= 10'b0;
      median_max_5_lpi_1_dfm_5 <= 3'b0;
      pixel_processing_pixel_processing_if_1_nor_itm_2 <= 1'b0;
      system_input_output_vld_sva_dfm_st_2 <= 1'b0;
      else_io_read_in_data_vld_rsc_svs_st_2 <= 1'b0;
      asn_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      buffer_slc_buffer_c_5_0_1_itm_2 <= 6'b0;
      buffer_acc_3_itm_2 <= 4'b0;
      buffer_acc_1_itm_2 <= 4'b0;
      else_io_read_in_data_vld_rsc_svs <= 1'b0;
      system_input_din_sva_1 <= 3'b0;
      buffer_t0_sva_1 <= 3'b0;
    end
    else begin
      out_data_rsci_ld <= and_dcpl_41 & asn_itm & (fsm_output[6]);
      in_data_rsci_ld <= and_159_cse;
      buffer_buf_buffer_buf_nor_itm_1 <= ~((buffer_buf_vinit_ndx_sva!=10'b0000000000));
      buffer_buf_acc_itm_2 <= nl_buffer_buf_acc_itm_2[9:0];
      median_max_5_lpi_1_dfm_5 <= MUX_v_3_2_2(median_max2_5_lpi_1_dfm_mx0, median_max2_6_lpi_1_dfm_mx0,
          and_131_nl);
      pixel_processing_pixel_processing_if_1_nor_itm_2 <= pixel_processing_pixel_processing_if_1_nor_itm;
      system_input_output_vld_sva_dfm_st_2 <= system_input_output_vld_sva_dfm_st_1;
      else_io_read_in_data_vld_rsc_svs_st_2 <= else_io_read_in_data_vld_rsc_svs_st_1;
      asn_itm_1 <= asn_itm;
      main_stage_0_2 <= ~ (fsm_output[2]);
      buffer_slc_buffer_c_5_0_1_itm_2 <= system_input_c_sva[5:0];
      buffer_acc_3_itm_2 <= nl_buffer_acc_3_itm_2[3:0];
      buffer_acc_1_itm_2 <= nl_buffer_acc_1_itm_2[3:0];
      else_io_read_in_data_vld_rsc_svs <= MUX_s_1_2_2(in_data_vld_rsci_d, else_io_read_in_data_vld_rsc_svs,
          or_tmp_49);
      system_input_din_sva_1 <= in_data_rsci_d;
      buffer_t0_sva_1 <= buffer_buf_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      buffer_buf_vinit_ndx_sva <= 10'b1001111111;
    end
    else if ( fsm_output[2] ) begin
      buffer_buf_vinit_ndx_sva <= buffer_buf_acc_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_7_sva <= 3'b0;
      system_input_window_6_sva <= 3'b0;
    end
    else if ( or_tmp_35 ) begin
      system_input_window_7_sva <= buffer_qr_1_lpi_1_dfm_mx0;
      system_input_window_6_sva <= buffer_qr_lpi_1_dfm_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_threshold_sva <= 3'b100;
    end
    else if ( and_12_itm & (fsm_output[5]) ) begin
      pixel_processing_threshold_sva <= mcu_data_rsci_q_d[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_r_sva <= 8'b0;
    end
    else if ( ~(or_dcpl_75 | (~((system_input_c_sva[8]) & (system_input_c_sva[5])
        & (system_input_c_sva[4]))) | (~((system_input_c_sva[3:1]==3'b111))) | or_dcpl_1
        | (~ (fsm_output[3]))) ) begin
      system_input_r_sva <= MUX_v_8_2_2(8'b00000000, (system_input_if_2_qelse_acc_nl),
          (system_input_if_2_system_input_if_2_nand_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_frame_sva <= 32'b1;
    end
    else if ( ~(and_dcpl_101 | (system_input_c_filter_sva[6]) | (system_input_c_filter_sva[7])
        | (~ (system_input_c_filter_sva[0])) | (~ (system_input_c_filter_sva[1]))
        | (~ (system_input_c_filter_sva[2])) | (~ (system_input_c_filter_sva[3]))
        | or_dcpl_87 | (~ (system_input_c_filter_sva[8])) | (~ in_data_vld_rsci_d)
        | (~ mcu_ready_sva) | (system_input_r_filter_sva[4]) | (~ (system_input_r_filter_sva[0]))
        | or_dcpl_81 | or_dcpl_80 | (~ (fsm_output[3]))) ) begin
      pixel_processing_frame_sva <= nl_pixel_processing_frame_sva[31:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_8_sva <= 3'b0;
    end
    else if ( and_cse & (fsm_output[4]) ) begin
      system_input_window_8_sva <= in_data_rsci_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_4_sva <= 3'b0;
    end
    else if ( ~ or_62_cse ) begin
      system_input_window_4_sva <= system_input_window_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_c_filter_sva <= 9'b0;
    end
    else if ( ~ or_62_cse ) begin
      system_input_c_filter_sva <= system_input_c_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_3_sva <= 3'b0;
    end
    else if ( ~ or_62_cse ) begin
      system_input_window_3_sva <= system_input_window_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_window_5_sva <= 3'b0;
    end
    else if ( ~ or_62_cse ) begin
      system_input_window_5_sva <= system_input_window_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_r_filter_sva <= 8'b0;
    end
    else if ( ~(and_dcpl_101 | (system_input_c_filter_sva[6]) | (system_input_c_filter_sva[7])
        | (~ (system_input_c_filter_sva[0])) | (~ (system_input_c_filter_sva[1]))
        | (~ (system_input_c_filter_sva[2])) | (~ (system_input_c_filter_sva[3]))
        | or_dcpl_87 | (~ (system_input_c_filter_sva[8])) | or_dcpl_1 | (~ (fsm_output[3])))
        ) begin
      system_input_r_filter_sva <= MUX_v_8_2_2(8'b00000000, (system_input_if_1_qelse_acc_nl),
          (clip_window_not_6_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_c_sva <= 9'b0;
    end
    else if ( ~ or_62_cse ) begin
      system_input_c_sva <= MUX_v_9_2_2(9'b000000000, (system_input_else_2_acc_nl),
          (system_input_system_input_nand_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_output_vld_sva <= 1'b0;
    end
    else if ( reg_system_input_system_input_output_vld_and_cse ) begin
      system_input_output_vld_sva <= system_input_output_vld_sva_dfm_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      mcu_ready_sva <= 1'b0;
    end
    else if ( fsm_output[5] ) begin
      mcu_ready_sva <= if_if_if_and_tmp | mcu_ready_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_pixel_processing_if_1_nor_itm <= 1'b0;
      system_input_output_vld_sva_dfm_st_1 <= 1'b0;
      else_io_read_in_data_vld_rsc_svs_st_1 <= 1'b0;
    end
    else if ( reg_pixel_processing_pixel_processing_if_1_pixel_processing_if_1_and_cse
        ) begin
      pixel_processing_pixel_processing_if_1_nor_itm <= ~((pixel_processing_mod10_acc_3_tmp!=3'b000)
          | (pixel_processing_frame_sva[0]));
      system_input_output_vld_sva_dfm_st_1 <= system_input_output_vld_sva_dfm_mx1w0;
      else_io_read_in_data_vld_rsc_svs_st_1 <= in_data_vld_rsci_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_asn_itm <= 3'b0;
      L2_5_L1a_4_slc_3_itm <= 1'b0;
      L2_5_L1a_3_slc_3_itm <= 1'b0;
    end
    else if ( pixel_processing_and_cse ) begin
      pixel_processing_asn_itm <= pixel_processing_threshold_sva;
      L2_5_L1a_4_slc_3_itm <= z_out_3;
      L2_5_L1a_3_slc_3_itm <= readslicef_4_1_3((L1a_if_acc_15_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_7_lpi_1_dfm <= 3'b0;
    end
    else if ( (mcu_ready_sva & z_out_3_3 & (fsm_output[5])) | and_133_rgt ) begin
      median_max_7_lpi_1_dfm <= MUX_v_3_2_2(median_max2_7_lpi_1_dfm_mx0, median_max2_8_lpi_1_dfm_mx0,
          and_133_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_6_lpi_1_dfm <= 3'b0;
      median_max_5_3_lpi_1_dfm <= 3'b0;
    end
    else if ( reg_median_median_max_or_2_cse ) begin
      median_max_6_lpi_1_dfm <= MUX_v_3_2_2(median_max2_6_3_lpi_1_dfm_mx0, L1b_asn_5_mx1w1,
          median_max_and_7_rgt);
      median_max_5_3_lpi_1_dfm <= MUX_v_3_2_2(L1b_asn_5_mx1w1, median_max2_6_3_lpi_1_dfm_mx0,
          median_max_and_7_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_4_1_lpi_1_dfm <= 3'b0;
    end
    else if ( (mcu_ready_sva & L1b_if_acc_10_itm_3 & (fsm_output[5])) | and_137_rgt
        ) begin
      median_max_4_1_lpi_1_dfm <= MUX_v_3_2_2(median_max2_4_lpi_1_dfm_mx0, median_max_2_lpi_1_dfm_mx0,
          and_137_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      buffer_sel_1_sva <= 1'b0;
    end
    else if ( reg_system_input_system_input_output_vld_and_cse | (fsm_output[2])
        ) begin
      buffer_sel_1_sva <= buffer_sel_1_sva_dfm_mx0 | (~(mcu_ready_sva & (fsm_output[3])));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      asn_itm <= 1'b0;
    end
    else if ( (fsm_output[2]) | (fsm_output[6]) ) begin
      asn_itm <= mcu_ready_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      clip_window_ac_int_cctor_2_sva_1 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      clip_window_ac_int_cctor_2_sva_1 <= and_146_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_if_2_asn_itm <= 32'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      pixel_processing_if_2_asn_itm <= pixel_processing_frame_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      pixel_processing_if_2_land_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      pixel_processing_if_2_land_lpi_1_dfm_1 <= pixel_processing_if_2_land_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_land_1_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      system_input_land_1_lpi_1_dfm_1 <= system_input_land_1_lpi_1_dfm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max2_1_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max2_1_lpi_1_dfm <= MUX_v_3_2_2(median_max2_0_lpi_1_dfm_1_mx0, median_max_1_2_lpi_1_dfm_mx0,
          median_max2_and_5_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_2_2_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max_2_2_lpi_1_dfm <= MUX_v_3_2_2(L1b_asn_44_mx0w1, median_max2_2_2_lpi_1_dfm_mx0,
          median_max_and_3_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max2_3_2_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max2_3_2_lpi_1_dfm <= MUX_v_3_2_2(median_max_2_1_lpi_1_dfm_mx0, median_max_3_1_lpi_1_dfm_mx0,
          median_max2_and_3_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max_4_2_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max_4_2_lpi_1_dfm <= MUX_v_3_2_2(median_max2_3_1_lpi_1_dfm_mx0, median_max2_4_1_lpi_1_dfm_mx0,
          median_max_and_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      median_max2_5_1_lpi_1_dfm <= 3'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      median_max2_5_1_lpi_1_dfm <= MUX_v_3_2_2(system_input_window_8_sva, system_input_window_7_sva,
          median_max2_median_max2_nor_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      clip_window_unequal_tmp_2 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      clip_window_unequal_tmp_2 <= (system_input_r_filter_sva!=8'b00000000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      clip_window_clip_window_and_1_cse_sva_1 <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      clip_window_clip_window_and_1_cse_sva_1 <= clip_window_clip_window_and_1_cse_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      system_input_output_vld_sva_dfm <= 1'b0;
    end
    else if ( ~ or_tmp_49 ) begin
      system_input_output_vld_sva_dfm <= system_input_output_vld_sva_dfm_mx1w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      buffer_sel_1_sva_dfm <= 1'b0;
    end
    else if ( ~ (fsm_output[4]) ) begin
      buffer_sel_1_sva_dfm <= buffer_sel_1_sva_dfm_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      and_cse <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      and_cse <= and_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      and_12_itm <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      and_12_itm <= pixel_processing_if_2_land_lpi_1_dfm & system_input_land_1_lpi_1_dfm
          & system_input_output_vld_sva_dfm_mx1w0 & in_data_vld_rsci_d & mcu_ready_sva;
    end
  end
  assign nl_buffer_buf_acc_itm_2  = buffer_buf_vinit_ndx_sva + 10'b1111111111;
  assign and_131_nl = and_dcpl_41 & (~ z_out_3_3);
  assign nl_buffer_acc_3_itm_2  = conv_u2u_3_4({buffer_sel_1_sva_dfm_mx0 , 1'b0 ,
      buffer_sel_1_sva_dfm_mx0}) + conv_u2u_3_4(system_input_c_sva[8:6]);
  assign nl_buffer_acc_1_itm_2  = conv_u2u_3_4(system_input_c_sva[8:6]) + 4'b101;
  assign nl_system_input_if_2_qelse_acc_nl = system_input_r_sva + 8'b1;
  assign system_input_if_2_qelse_acc_nl = nl_system_input_if_2_qelse_acc_nl[7:0];
  assign system_input_if_2_system_input_if_2_nand_nl = ~((system_input_r_sva==8'b11101111));
  assign nl_pixel_processing_frame_sva  = pixel_processing_frame_sva + 32'b1;
  assign nl_system_input_if_1_qelse_acc_nl = system_input_r_filter_sva + 8'b1;
  assign system_input_if_1_qelse_acc_nl = nl_system_input_if_1_qelse_acc_nl[7:0];
  assign clip_window_not_6_nl = ~ and_146_cse;
  assign nl_system_input_else_2_acc_nl = system_input_c_sva + 9'b1;
  assign system_input_else_2_acc_nl = nl_system_input_else_2_acc_nl[8:0];
  assign system_input_system_input_nand_nl = ~((system_input_c_sva==9'b100111111));
  assign L1b_mux_2_nl = MUX_v_3_2_2(median_max_2_lpi_1_dfm_mx0, median_max2_4_lpi_1_dfm_mx0,
      L1b_if_acc_10_itm_3);
  assign L1b_mux_3_nl = MUX_v_3_2_2(median_max2_6_3_lpi_1_dfm_mx0, L1b_asn_5_mx1w1,
      L1b_if_acc_11_itm_3);
  assign nl_L1a_if_acc_15_nl = ({1'b1 , (L1b_mux_2_nl)}) + conv_u2u_3_4(~ (L1b_mux_3_nl))
      + 4'b1;
  assign L1a_if_acc_15_nl = nl_L1a_if_acc_15_nl[3:0];
  assign median_max2_and_5_nl = z_out_3 & (~ (fsm_output[4]));
  assign median_max_and_3_nl = z_out_3_3 & (~ (fsm_output[4]));
  assign median_max2_and_3_nl = z_out_2_3 & (~ (fsm_output[4]));
  assign median_max_and_1_nl = z_out_4_3 & (~ (fsm_output[4]));
  assign median_max2_median_max2_nor_nl = ~((~(and_146_cse | (~ z_out_5_3))) | (fsm_output[4]));
  assign thresholding_if_and_2_nl = (~ L1b_if_acc_11_itm_3) & (fsm_output[5]);
  assign thresholding_if_and_3_nl = L1b_if_acc_11_itm_3 & (fsm_output[5]);
  assign thresholding_if_mux1h_3_nl = MUX1HOT_v_3_4_2((~ pixel_processing_asn_itm),
      median_max2_0_lpi_1_dfm_1_mx0, L1b_asn_5_mx1w1, median_max2_6_3_lpi_1_dfm_mx0,
      {(fsm_output[6]) , (fsm_output[3]) , (thresholding_if_and_2_nl) , (thresholding_if_and_3_nl)});
  assign L1b_mux_30_nl = MUX_v_3_2_2(median_max2_8_lpi_1_dfm_mx0, median_max2_7_lpi_1_dfm_mx0,
      z_out_3_3);
  assign thresholding_if_mux1h_4_nl = MUX1HOT_v_3_3_2(median_max_5_lpi_1_dfm_mx0,
      (~ median_max_1_2_lpi_1_dfm_mx0), (~ (L1b_mux_30_nl)), {(fsm_output[6]) , (fsm_output[3])
      , (fsm_output[5])});
  assign nl_acc_nl = ({1'b1 , (thresholding_if_mux1h_3_nl) , 1'b1}) + conv_u2u_4_5({(thresholding_if_mux1h_4_nl)
      , 1'b1});
  assign acc_nl = nl_acc_nl[4:0];
  assign z_out_3 = readslicef_5_1_4((acc_nl));
  assign L1a_if_mux_19_nl = MUX_v_3_2_2(pixel_processing_window_2_lpi_1_dfm_mx0,
      median_max_4_2_lpi_1_dfm, fsm_output[5]);
  assign L1a_if_mux_20_nl = MUX_v_3_2_2((~ clip_window_qr_3_lpi_1_dfm_mx0), (~ median_max_5_2_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_1_nl = ({1'b1 , (L1a_if_mux_19_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux_20_nl)
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[4:0];
  assign z_out_1_3 = readslicef_5_1_4((acc_1_nl));
  assign L1a_if_mux_21_nl = MUX_v_3_2_2(median_max_8_lpi_1_dfm_mx0, median_max_2_1_lpi_1_dfm_mx0,
      fsm_output[3]);
  assign L1a_if_mux_22_nl = MUX_v_3_2_2((~ median_max2_9_lpi_1_dfm_1_mx0), (~ median_max_3_1_lpi_1_dfm_mx0),
      fsm_output[3]);
  assign nl_acc_2_nl = ({1'b1 , (L1a_if_mux_21_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux_22_nl)
      , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[4:0];
  assign z_out_2_3 = readslicef_5_1_4((acc_2_nl));
  assign L1b_if_mux1h_3_nl = MUX1HOT_v_3_3_2(median_max2_5_lpi_1_dfm_mx0, median_max2_7_lpi_1_dfm_mx0,
      L1b_asn_44_mx0w1, {(fsm_output[6]) , (fsm_output[5]) , (fsm_output[3])});
  assign L1b_if_mux1h_4_nl = MUX1HOT_v_3_3_2((~ median_max2_6_lpi_1_dfm_mx0), (~
      median_max2_8_lpi_1_dfm_mx0), (~ median_max2_2_2_lpi_1_dfm_mx0), {(fsm_output[6])
      , (fsm_output[5]) , (fsm_output[3])});
  assign nl_acc_3_nl = ({1'b1 , (L1b_if_mux1h_3_nl) , 1'b1}) + conv_u2u_4_5({(L1b_if_mux1h_4_nl)
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[4:0];
  assign z_out_3_3 = readslicef_5_1_4((acc_3_nl));
  assign L1b_if_mux_6_nl = MUX_v_3_2_2(median_max2_3_1_lpi_1_dfm_mx0, median_max2_3_2_lpi_1_dfm,
      fsm_output[5]);
  assign L1b_if_mux_7_nl = MUX_v_3_2_2((~ median_max2_4_1_lpi_1_dfm_mx0), (~ median_max2_4_2_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_4_nl = ({1'b1 , (L1b_if_mux_6_nl) , 1'b1}) + conv_u2u_4_5({(L1b_if_mux_7_nl)
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[4:0];
  assign z_out_4_3 = readslicef_5_1_4((acc_4_nl));
  assign L1a_if_mux_23_nl = MUX_v_3_2_2(system_input_window_7_sva, median_max2_7_1_lpi_1_dfm_mx0,
      fsm_output[5]);
  assign clip_window_mux_8_nl = MUX_v_3_2_2(system_input_window_8_sva, system_input_window_7_sva,
      and_146_cse);
  assign L1a_if_mux_24_nl = MUX_v_3_2_2((~ (clip_window_mux_8_nl)), (~ pixel_processing_window_8_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_5_nl = ({1'b1 , (L1a_if_mux_23_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux_24_nl)
      , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[4:0];
  assign z_out_5_3 = readslicef_5_1_4((acc_5_nl));
  assign L1a_if_mux_25_nl = MUX_v_3_2_2(median_max2_0_lpi_1_dfm_mx0, L1a_asn_13_mx0w1,
      fsm_output[5]);
  assign L1a_if_mux_26_nl = MUX_v_3_2_2((~ median_max_1_1_lpi_1_dfm_mx0), (~ median_max_7_2_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_6_nl = ({1'b1 , (L1a_if_mux_25_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux_26_nl)
      , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[4:0];
  assign z_out_6_3 = readslicef_5_1_4((acc_6_nl));
  assign L1b_if_mux_8_nl = MUX_v_3_2_2(median_max2_1_1_lpi_1_dfm_mx0, median_max2_7_2_lpi_1_dfm_mx0,
      fsm_output[5]);
  assign L1b_if_mux_9_nl = MUX_v_3_2_2((~ median_max2_2_1_lpi_1_dfm_mx0), (~ median_max2_8_2_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_7_nl = ({1'b1 , (L1b_if_mux_8_nl) , 1'b1}) + conv_u2u_4_5({(L1b_if_mux_9_nl)
      , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[4:0];
  assign z_out_7_3 = readslicef_5_1_4((acc_7_nl));
  assign L1a_if_mux_27_nl = MUX_v_3_2_2(pixel_processing_window_0_lpi_1_dfm_mx0,
      median_max_8_1_lpi_1_dfm_mx0, fsm_output[5]);
  assign L1a_if_mux_28_nl = MUX_v_3_2_2((~ clip_window_qr_lpi_1_dfm_mx0), (~ median_max2_9_lpi_1_dfm_mx0),
      fsm_output[5]);
  assign nl_acc_8_nl = ({1'b1 , (L1a_if_mux_27_nl) , 1'b1}) + conv_u2u_4_5({(L1a_if_mux_28_nl)
      , 1'b1});
  assign acc_8_nl = nl_acc_8_nl[4:0];
  assign z_out_8_3 = readslicef_5_1_4((acc_8_nl));

  function [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function  [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function  [3:0] conv_s2s_2_4 ;
    input [1:0]  vector ;
  begin
    conv_s2s_2_4 = {{2{vector[1]}}, vector};
  end
  endfunction


  function  [2:0] conv_s2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_3 = {vector[1], vector};
  end
  endfunction


  function  [3:0] conv_s2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2u_3_4 = {vector[2], vector};
  end
  endfunction


  function  [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction


  function  [3:0] conv_u2s_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2s_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function  [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function  [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction


  function  [5:0] conv_u2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    filter
// ------------------------------------------------------------------


module filter (
  clk, rst, in_data_rsc_z, in_data_rsc_lz, in_data_vld_rsc_z, out_data_rsc_z, out_data_rsc_lz,
      mcu_data_rsc_adr, mcu_data_rsc_q, mcu_data_rsc_d, mcu_data_rsc_we
);
  input clk;
  input rst;
  input [2:0] in_data_rsc_z;
  output in_data_rsc_lz;
  input in_data_vld_rsc_z;
  output [2:0] out_data_rsc_z;
  output out_data_rsc_lz;
  output [8:0] mcu_data_rsc_adr;
  input [31:0] mcu_data_rsc_q;
  output [31:0] mcu_data_rsc_d;
  output mcu_data_rsc_we;


  // Interconnect Declarations
  wire [8:0] mcu_data_rsci_adr_d;
  wire [31:0] mcu_data_rsci_d_d;
  wire mcu_data_rsci_we_d;
  wire [31:0] mcu_data_rsci_q_d;
  wire mcu_data_rsci_ram_rw_A_internal_RMASK_B_d;
  wire [9:0] buffer_buf_rsci_radr_d;
  wire [9:0] buffer_buf_rsci_wadr_d;
  wire [2:0] buffer_buf_rsci_d_d;
  wire buffer_buf_rsci_we_d;
  wire buffer_buf_rsci_re_d;
  wire [2:0] buffer_buf_rsci_q_d;
  wire buffer_buf_rsc_we;
  wire [2:0] buffer_buf_rsc_d;
  wire [9:0] buffer_buf_rsc_wadr;
  wire buffer_buf_rsc_re;
  wire [2:0] buffer_buf_rsc_q;
  wire [9:0] buffer_buf_rsc_radr;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.data_width(32'sd3),
  .addr_width(32'sd10),
  .depth(32'sd640)) buffer_buf_rsc_comp (
      .radr(buffer_buf_rsc_radr),
      .wadr(buffer_buf_rsc_wadr),
      .d(buffer_buf_rsc_d),
      .we(buffer_buf_rsc_we),
      .re(buffer_buf_rsc_re),
      .clk(clk),
      .q(buffer_buf_rsc_q)
    );
  Xilinx_RAMS_BLOCK_SPRAM_RBW_rwport_32_9_512_4_gen mcu_data_rsci (
      .we(mcu_data_rsc_we),
      .d(mcu_data_rsc_d),
      .q(mcu_data_rsc_q),
      .adr(mcu_data_rsc_adr),
      .adr_d(mcu_data_rsci_adr_d),
      .d_d(mcu_data_rsci_d_d),
      .we_d(mcu_data_rsci_we_d),
      .q_d(mcu_data_rsci_q_d),
      .ram_rw_A_internal_RMASK_B_d(mcu_data_rsci_ram_rw_A_internal_RMASK_B_d)
    );
  Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_10_640_7_gen buffer_buf_rsci (
      .we(buffer_buf_rsc_we),
      .d(buffer_buf_rsc_d),
      .wadr(buffer_buf_rsc_wadr),
      .re(buffer_buf_rsc_re),
      .q(buffer_buf_rsc_q),
      .radr(buffer_buf_rsc_radr),
      .radr_d(buffer_buf_rsci_radr_d),
      .wadr_d(buffer_buf_rsci_wadr_d),
      .d_d(buffer_buf_rsci_d_d),
      .we_d(buffer_buf_rsci_we_d),
      .re_d(buffer_buf_rsci_re_d),
      .q_d(buffer_buf_rsci_q_d)
    );
  filter_core filter_core_inst (
      .clk(clk),
      .rst(rst),
      .in_data_rsc_z(in_data_rsc_z),
      .in_data_rsc_lz(in_data_rsc_lz),
      .in_data_vld_rsc_z(in_data_vld_rsc_z),
      .out_data_rsc_z(out_data_rsc_z),
      .out_data_rsc_lz(out_data_rsc_lz),
      .mcu_data_rsci_adr_d(mcu_data_rsci_adr_d),
      .mcu_data_rsci_d_d(mcu_data_rsci_d_d),
      .mcu_data_rsci_we_d(mcu_data_rsci_we_d),
      .mcu_data_rsci_q_d(mcu_data_rsci_q_d),
      .mcu_data_rsci_ram_rw_A_internal_RMASK_B_d(mcu_data_rsci_ram_rw_A_internal_RMASK_B_d),
      .buffer_buf_rsci_radr_d(buffer_buf_rsci_radr_d),
      .buffer_buf_rsci_wadr_d(buffer_buf_rsci_wadr_d),
      .buffer_buf_rsci_d_d(buffer_buf_rsci_d_d),
      .buffer_buf_rsci_we_d(buffer_buf_rsci_we_d),
      .buffer_buf_rsci_re_d(buffer_buf_rsci_re_d),
      .buffer_buf_rsci_q_d(buffer_buf_rsci_q_d)
    );
endmodule



