
//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_in_wire_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


`ifdef mgc_in_wire_v1
`else
`define mgc_in_wire_v1
module mgc_in_wire_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule
`endif


//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/siflibs/mgc_out_stdreg_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

`ifdef mgc_out_stdreg_v1
`else
`define mgc_out_stdreg_v1
module mgc_out_stdreg_v1 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule
`endif




//------> C:/PROGRA~1/MENTOR~1/CATAPU~1.0C/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW.v 
// Block 1R1W Read Before Write RAM with common clock
`ifdef BLOCK_1R1W_RBW
`else
`define BLOCK_1R1W_RBW
module BLOCK_1R1W_RBW
#(
parameter data_width = 8,
parameter addr_width = 7,
parameter depth = 128
)(
	radr, wadr, d, we, re, clk, q
);

	input [addr_width-1:0] radr;
	input [addr_width-1:0] wadr;
	input [data_width-1:0] d;
	input we;
	input re;
	input clk;
	output[data_width-1:0] q;

	reg [data_width-1:0] q;

	(* ram_style = "block" *)
	reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block_ram"
	//pragma attribute mem block_ram true
		
	always @(posedge clk) begin
		if (we) begin
			mem[wadr] <= d; // Write port
		end
		if (re) begin
			q <= mem[radr] ; // read port
		end
	end

endmodule
`endif

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0c/745553 Production Release
//  HLS Date:       Wed Oct 11 16:38:17 PDT 2017
// 
//  Generated by:   Fitkit@DESKTOP-NJUNEBJ
//  Generated date: Tue Oct 31 12:27:49 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_11_1280_8_gen
// ------------------------------------------------------------------


`ifdef Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_11_1280_8_gen
`else
`define Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_11_1280_8_gen
module Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_11_1280_8_gen (
  we, d, wadr, re, q, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d
);
  output we;
  output [2:0] d;
  output [10:0] wadr;
  output re;
  input [2:0] q;
  output [10:0] radr;
  input [10:0] radr_d;
  input [10:0] wadr_d;
  input [2:0] d_d;
  input we_d;
  input re_d;
  output [2:0] q_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (we_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign re = (re_d);
  assign q_d = q;
  assign radr = (radr_d);
endmodule
`endif

// ------------------------------------------------------------------
//  Design Unit:    video_buf_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


`ifdef video_buf_core_core_fsm
`else
`define video_buf_core_core_fsm
module video_buf_core_core_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for video_buf_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : video_buf_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= core_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule
`endif

// ------------------------------------------------------------------
//  Design Unit:    video_buf_core
// ------------------------------------------------------------------


`ifdef video_buf_core
`else
`define video_buf_core
module video_buf_core (
  clk, rst, in_data_rsc_z, in_data_vld_rsc_z, vga_row_rsc_z, vga_col_rsc_z, out_data_rsc_z,
      vga_enable_rsc_z, gen_pause_rsc_z, buffer_rsci_radr_d, buffer_rsci_wadr_d,
      buffer_rsci_d_d, buffer_rsci_we_d, buffer_rsci_re_d, buffer_rsci_q_d
);
  input clk;
  input rst;
  input [2:0] in_data_rsc_z;
  input in_data_vld_rsc_z;
  input [9:0] vga_row_rsc_z;
  input [9:0] vga_col_rsc_z;
  output [2:0] out_data_rsc_z;
  output vga_enable_rsc_z;
  output gen_pause_rsc_z;
  output [10:0] buffer_rsci_radr_d;
  output [10:0] buffer_rsci_wadr_d;
  output [2:0] buffer_rsci_d_d;
  output buffer_rsci_we_d;
  output buffer_rsci_re_d;
  input [2:0] buffer_rsci_q_d;


  // Interconnect Declarations
  wire [2:0] in_data_rsci_d;
  wire in_data_vld_rsci_d;
  wire [9:0] vga_row_rsci_d;
  wire [9:0] vga_col_rsci_d;
  reg [2:0] out_data_rsci_d;
  reg vga_enable_rsci_d;
  reg gen_pause_rsci_d;
  wire [1:0] fsm_output;
  wire or_tmp_1;
  reg [1:0] row_in_sva;
  wire [2:0] nl_row_in_sva;
  reg [9:0] col_in_sva;
  reg vga_enable_int_sva_dfm_2;
  reg and_itm_2;
  reg reg_buffer_rsci_re_d_cse;

  wire[9:0] if_2_else_acc_nl;
  wire[10:0] nl_if_2_else_acc_nl;
  wire[0:0] if_2_if_2_nand_nl;
  wire[4:0] and_21_nl;
  wire[4:0] acc_3_nl;
  wire[5:0] nl_acc_3_nl;
  wire[5:0] vga_col_vga_col_and_nl;
  wire[4:0] if_2_if_2_and_2_nl;
  wire[4:0] if_2_acc_nl;
  wire[5:0] nl_if_2_acc_nl;
  wire[5:0] if_2_if_2_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire_v1 #(.rscid(32'sd1),
  .width(32'sd3)) in_data_rsci (
      .d(in_data_rsci_d),
      .z(in_data_rsc_z)
    );
  mgc_in_wire_v1 #(.rscid(32'sd2),
  .width(32'sd1)) in_data_vld_rsci (
      .d(in_data_vld_rsci_d),
      .z(in_data_vld_rsc_z)
    );
  mgc_in_wire_v1 #(.rscid(32'sd3),
  .width(32'sd10)) vga_row_rsci (
      .d(vga_row_rsci_d),
      .z(vga_row_rsc_z)
    );
  mgc_in_wire_v1 #(.rscid(32'sd4),
  .width(32'sd10)) vga_col_rsci (
      .d(vga_col_rsci_d),
      .z(vga_col_rsc_z)
    );
  mgc_out_stdreg_v1 #(.rscid(32'sd5),
  .width(32'sd3)) out_data_rsci (
      .d(out_data_rsci_d),
      .z(out_data_rsc_z)
    );
  mgc_out_stdreg_v1 #(.rscid(32'sd6),
  .width(32'sd1)) vga_enable_rsci (
      .d(vga_enable_rsci_d),
      .z(vga_enable_rsc_z)
    );
  mgc_out_stdreg_v1 #(.rscid(32'sd7),
  .width(32'sd1)) gen_pause_rsci (
      .d(gen_pause_rsci_d),
      .z(gen_pause_rsc_z)
    );
  video_buf_core_core_fsm video_buf_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign or_tmp_1 = in_data_vld_rsci_d & (fsm_output[1]);
  assign nl_acc_3_nl = conv_u2u_3_5(vga_col_rsci_d[9:7]) + conv_u2u_4_5({(vga_row_rsci_d[2:1])
      , (vga_row_rsci_d[2:1])});
  assign acc_3_nl = nl_acc_3_nl[4:0];
  assign and_21_nl = MUX_v_5_2_2(5'b00000, (acc_3_nl), (fsm_output[1]));
  assign vga_col_vga_col_and_nl = MUX_v_6_2_2(6'b000000, (vga_col_rsci_d[6:1]), (fsm_output[1]));
  assign buffer_rsci_radr_d = {(and_21_nl) , (vga_col_vga_col_and_nl)};
  assign nl_if_2_acc_nl = conv_u2u_4_5(col_in_sva[9:6]) + conv_u2u_4_5({row_in_sva
      , row_in_sva});
  assign if_2_acc_nl = nl_if_2_acc_nl[4:0];
  assign if_2_if_2_and_2_nl = MUX_v_5_2_2(5'b00000, (if_2_acc_nl), or_tmp_1);
  assign if_2_if_2_and_1_nl = MUX_v_6_2_2(6'b000000, (col_in_sva[5:0]), or_tmp_1);
  assign buffer_rsci_wadr_d = {(if_2_if_2_and_2_nl) , (if_2_if_2_and_1_nl)};
  assign buffer_rsci_d_d = MUX_v_3_2_2(3'b000, in_data_rsci_d, or_tmp_1);
  assign buffer_rsci_we_d = or_tmp_1;
  assign buffer_rsci_re_d = fsm_output[1];
  always @(posedge clk) begin
    if ( rst ) begin
      gen_pause_rsci_d <= 1'b0;
      vga_enable_rsci_d <= 1'b0;
      out_data_rsci_d <= 3'b0;
    end
    else if ( reg_buffer_rsci_re_d_cse ) begin
      gen_pause_rsci_d <= and_itm_2;
      vga_enable_rsci_d <= vga_enable_int_sva_dfm_2;
      out_data_rsci_d <= buffer_rsci_q_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_buffer_rsci_re_d_cse <= 1'b0;
      and_itm_2 <= 1'b0;
      vga_enable_int_sva_dfm_2 <= 1'b0;
    end
    else begin
      reg_buffer_rsci_re_d_cse <= fsm_output[1];
      and_itm_2 <= (~(((~ (vga_row_rsci_d[1])) | (row_in_sva[0])) ^ (vga_row_rsci_d[2])
          ^ (row_in_sva[1]))) & ((vga_row_rsci_d[1]) ^ (row_in_sva[0]));
      vga_enable_int_sva_dfm_2 <= (vga_enable_int_sva_dfm_2 & reg_buffer_rsci_re_d_cse)
          | ((row_in_sva==2'b10));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      col_in_sva <= 10'b0;
    end
    else if ( ~((~ in_data_vld_rsci_d) | (fsm_output[0])) ) begin
      col_in_sva <= MUX_v_10_2_2(10'b0000000000, (if_2_else_acc_nl), (if_2_if_2_nand_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      row_in_sva <= 2'b0;
    end
    else if ( ~((~ in_data_vld_rsci_d) | (col_in_sva!=10'b0100111111)) ) begin
      row_in_sva <= nl_row_in_sva[1:0];
    end
  end
  assign nl_if_2_else_acc_nl = col_in_sva + 10'b1;
  assign if_2_else_acc_nl = nl_if_2_else_acc_nl[9:0];
  assign if_2_if_2_nand_nl = ~((col_in_sva==10'b0100111111));
  assign nl_row_in_sva  = row_in_sva + 2'b1;

  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function  [4:0] conv_u2u_3_5 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_5 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [4:0] conv_u2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction

endmodule
`endif

// ------------------------------------------------------------------
//  Design Unit:    video_buf
// ------------------------------------------------------------------


`ifdef video_buf
`else
`define video_buf
module video_buf (
  clk, rst, in_data_rsc_z, in_data_vld_rsc_z, vga_row_rsc_z, vga_col_rsc_z, out_data_rsc_z,
      vga_enable_rsc_z, gen_pause_rsc_z
);
  input clk;
  input rst;
  input [2:0] in_data_rsc_z;
  input in_data_vld_rsc_z;
  input [9:0] vga_row_rsc_z;
  input [9:0] vga_col_rsc_z;
  output [2:0] out_data_rsc_z;
  output vga_enable_rsc_z;
  output gen_pause_rsc_z;


  // Interconnect Declarations
  wire [10:0] buffer_rsci_radr_d;
  wire [10:0] buffer_rsci_wadr_d;
  wire [2:0] buffer_rsci_d_d;
  wire buffer_rsci_we_d;
  wire buffer_rsci_re_d;
  wire [2:0] buffer_rsci_q_d;
  wire buffer_rsc_we;
  wire [2:0] buffer_rsc_d;
  wire [10:0] buffer_rsc_wadr;
  wire buffer_rsc_re;
  wire [2:0] buffer_rsc_q;
  wire [10:0] buffer_rsc_radr;


  // Interconnect Declarations for Component Instantiations 
  BLOCK_1R1W_RBW #(.data_width(32'sd3),
  .addr_width(32'sd11),
  .depth(32'sd1280)) buffer_rsc_comp (
      .radr(buffer_rsc_radr),
      .wadr(buffer_rsc_wadr),
      .d(buffer_rsc_d),
      .we(buffer_rsc_we),
      .re(buffer_rsc_re),
      .clk(clk),
      .q(buffer_rsc_q)
    );
  Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_3_11_1280_8_gen buffer_rsci (
      .we(buffer_rsc_we),
      .d(buffer_rsc_d),
      .wadr(buffer_rsc_wadr),
      .re(buffer_rsc_re),
      .q(buffer_rsc_q),
      .radr(buffer_rsc_radr),
      .radr_d(buffer_rsci_radr_d),
      .wadr_d(buffer_rsci_wadr_d),
      .d_d(buffer_rsci_d_d),
      .we_d(buffer_rsci_we_d),
      .re_d(buffer_rsci_re_d),
      .q_d(buffer_rsci_q_d)
    );
  video_buf_core video_buf_core_inst (
      .clk(clk),
      .rst(rst),
      .in_data_rsc_z(in_data_rsc_z),
      .in_data_vld_rsc_z(in_data_vld_rsc_z),
      .vga_row_rsc_z(vga_row_rsc_z),
      .vga_col_rsc_z(vga_col_rsc_z),
      .out_data_rsc_z(out_data_rsc_z),
      .vga_enable_rsc_z(vga_enable_rsc_z),
      .gen_pause_rsc_z(gen_pause_rsc_z),
      .buffer_rsci_radr_d(buffer_rsci_radr_d),
      .buffer_rsci_wadr_d(buffer_rsci_wadr_d),
      .buffer_rsci_d_d(buffer_rsci_d_d),
      .buffer_rsci_we_d(buffer_rsci_we_d),
      .buffer_rsci_re_d(buffer_rsci_re_d),
      .buffer_rsci_q_d(buffer_rsci_q_d)
    );
endmodule
`endif



